module LUT1(
    input[4:0] addr,
    output logic[9:0] Target
	);

always_comb 
  case(addr)		   
	5'b00000:   Target =  10'b0000001011; //lut[0] = 11
	5'b00001:   Target =  10'b0010101001; //lut[1] = 169
	5'b00010:   Target =  10'b0100101110; //lut[2] = 302
	5'b00011:   Target =  10'b0100110001; //lut[3] = 305
	5'b00100:   Target =  10'b0100111010; //lut[4] = 314
	5'b00101:   Target =  10'b0100111101; //lut[5] = 317
	5'b00110:   Target =  10'b0101111101; //lut[6] = 381
	5'b00111:   Target =  10'b0110000010; //lut[7] = 386
	5'b01000:   Target =  10'b0110001000; //lut[8] = 392
	5'b01001:   Target =  10'b0110001111; //lut[9] = 399
	5'b01010:   Target =  10'b0110010111; //lut[10] = 407
	5'b01011:   Target =  10'b0110100000; //lut[11] = 416
	5'b01100:   Target =  10'b0111010010; //lut[12] = 446
	5'b01101:   Target =  10'b0111000100; //lut[13] = 452
	5'b01110:   Target =  10'b0111001011; //lut[14] = 459
	5'b01111:   Target =  10'b0111010011; //lut[15] = 467
	5'b10000:   Target =  10'b0111011100; //lut[16] = 476
	5'b10001:   Target =  10'b0111100110; //lut[17] = 486
	5'b10010:   Target =  10'b0111100110; //lut[18] = 486
	5'b10011:   Target =  10'b0111111101; //lut[19] = 509
	5'b10100:   Target =  10'b1000000001; //lut[20] = 513
	5'b10101:   Target =  10'b1000000110; //lut[21] = 518
	5'b10110:   Target =  10'b1000001011; //lut[22] = 523
	5'b10111:   Target =  10'b1000010000; //lut[23] = 528
	5'b11000:   Target =  10'b1000010101; //lut[24] = 533
	5'b11001:   Target =  10'b1000011000; //lut[25] = 536
	5'b11010:   Target =  10'b1000100000; //lut[26] = 544
	5'b11011:   Target =  10'b1000101000; //lut[26] = 552
	default: Target = 10'b0000000000;
  endcase
endmodule
